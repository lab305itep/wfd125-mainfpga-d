localparam VERSION = 32'h00030001;